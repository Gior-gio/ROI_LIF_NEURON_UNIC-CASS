** sch_path: /foss/designs/chipathon_2025/designs/ihp-sg13g2/edge_detector/xschem/edge_detector.sch
.subckt edge_detector IN OUT VDD VSS
*.PININFO VDD:B VSS:B IN:I OUT:O
xINV0 VDD I0 IN VSS gate_inv_L0d5
xINV1 VDD I1 I0 VSS gate_inv_L0d5
xINV2 VDD I2 I1 VSS gate_inv_L0d5
xINV3 VDD I3 I2 VSS gate_inv_L0d5
xINV4 VDD I4 I3 VSS gate_inv_L0d5
xAND IN VDD VSS OUT I4 gate_and
.ends

* expanding   symbol:  /foss/designs/chipathon_2025/designs/ihp-sg13g2/gate_inv_L0d5/xschem/gate_inv_L0d5.sym # of pins=4
** sym_path: /foss/designs/chipathon_2025/designs/ihp-sg13g2/gate_inv_L0d5/xschem/gate_inv_L0d5.sym
** sch_path: /foss/designs/chipathon_2025/designs/ihp-sg13g2/gate_inv_L0d5/xschem/gate_inv_L0d5.sch
.subckt gate_inv_L0d5 VDD B A VSS
*.PININFO B:O A:I VDD:B VSS:B
XMN B A VSS VSS sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XMP B A VDD VDD sg13_lv_pmos w=2u l=0.5u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/chipathon_2025/designs/ihp-sg13g2/gate_and/xschem/gate_and.sym # of pins=5
** sym_path: /foss/designs/chipathon_2025/designs/ihp-sg13g2/gate_and/xschem/gate_and.sym
** sch_path: /foss/designs/chipathon_2025/designs/ihp-sg13g2/gate_and/xschem/gate_and.sch
.subckt gate_and B VDD VSS OUT A
*.PININFO OUT:O A:I VDD:B VSS:B B:I
XMNB OUTN B NX VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMNA NX A VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMPB OUTN B VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XMPA OUTN A VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XMNI OUT OUTN VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMPI OUT OUTN VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
.ends

