* Extracted by KLayout with GF180MCU LVS runset on : 15/11/2025 23:55

.SUBCKT gate_or VSS B OUTN OUT A VDD
M$1 \$32 A VDD VDD pfet_03v3 L=0.28U W=12U AS=6.06P AD=5.16P PS=19.04U PD=15.44U
M$5 \$32 VDD VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$6 OUTN B \$32 VDD pfet_03v3 L=0.28U W=12U AS=5.16P AD=5.16P PS=15.44U
+ PD=15.44U
M$11 OUT OUTN VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=3.48P PS=7.72U
+ PD=11.32U
M$13 VSS VSS VSS VSS nfet_03v3 L=0.28U W=4U AS=2.02P AD=1.72P PS=9.04U PD=7.44U
M$14 OUTN A VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$18 OUTN VSS VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$19 VSS B OUTN VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$23 OUT OUTN VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=1.16P PS=3.72U PD=5.32U
.ENDS gate_or
