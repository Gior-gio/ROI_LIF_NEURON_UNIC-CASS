** sch_path: /foss/designs/chipathon_2025/designs/gf180/spike_generator/spike_generator.sch
.subckt spike_generator VDD Vcmp Vspk Vrst Ven VSS
*.PININFO Vcmp:B Ven:B Vrst:B Vspk:B VDD:B VSS:B
xOR Ven VDD VSS X VCMPB gate_or
xED VCMPB SPK_OUT VDD VSS edge_detector_TOP
xBUF2 VDD Vspk SPK_OUT VSS gate_buf_L0d28
x1 VDD VCMPB Vcmp VSS gate_inv_L0d28
xBUF1 VDD Vrst X VSS gate_buf_L0d28
.ends

* expanding   symbol:  gf180/gate_or/xschem/gate_or.sym # of pins=5
** sym_path: /foss/designs/chipathon_2025/designs/gf180/gate_or/xschem/gate_or.sym
** sch_path: /foss/designs/chipathon_2025/designs/gf180/gate_or/xschem/gate_or.sch
.subckt gate_or B VDD VSS OUT A
*.PININFO OUT:O A:I VDD:B VSS:B B:I
MNB OUTN B VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MPB OUTN B net1 VDD pfet_03v3 L=0.28u W=3u nf=1 m=4
MNA OUTN A VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MPA net1 A VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=4
MIN OUT OUTN VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MIP OUT OUTN VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
MPB1 net1 VDD VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
MNA1 OUTN VSS VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MNA2 VSS VSS VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=4
.ends


* expanding   symbol:  gf180/edge_detector/xschem/edge_detector_TOP.sym # of pins=4
** sym_path: /foss/designs/chipathon_2025/designs/gf180/edge_detector/xschem/edge_detector_TOP.sym
** sch_path: /foss/designs/chipathon_2025/designs/gf180/edge_detector/xschem/edge_detector_TOP.sch
.subckt edge_detector_TOP IN OUT VDD VSS
*.PININFO VDD:B VSS:B IN:I OUT:O
xAND IN VDD VSS OUT X[4] gate_and
xINV0 VDD X[0] IN VSS gate_inv_L0d5
xINV1 VDD X[1] X[0] VSS gate_inv_L0d5
xINV2 VDD X[2] X[1] VSS gate_inv_L0d5
xINV3 VDD X[3] X[2] VSS gate_inv_L0d5
xINV4 VDD X[4] X[3] VSS gate_inv_L0d5
.ends


* expanding   symbol:  gf180/gate_buf_L0d28/xschem/gate_buf_L0d28.sym # of pins=4
** sym_path: /foss/designs/chipathon_2025/designs/gf180/gate_buf_L0d28/xschem/gate_buf_L0d28.sym
** sch_path: /foss/designs/chipathon_2025/designs/gf180/gate_buf_L0d28/xschem/gate_buf_L0d28.sch
.subckt gate_buf_L0d28 VDD B A VSS
*.PININFO B:O A:I VDD:B VSS:B
MN1 net1 A VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MP1 net1 A VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
MN2 B net1 VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=6
MP2 B net1 VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=6
.ends


* expanding   symbol:  gf180/gate_inv_L0d28/xschem/gate_inv_L0d28.sym # of pins=4
** sym_path: /foss/designs/chipathon_2025/designs/gf180/gate_inv_L0d28/xschem/gate_inv_L0d28.sym
** sch_path: /foss/designs/chipathon_2025/designs/gf180/gate_inv_L0d28/xschem/gate_inv_L0d28.sch
.subckt gate_inv_L0d28 VDD B A VSS
*.PININFO B:O A:I VDD:B VSS:B
MN B A VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MP B A VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
.ends


* expanding   symbol:  gf180/gate_and/xschem/gate_and.sym # of pins=5
** sym_path: /foss/designs/chipathon_2025/designs/gf180/gate_and/xschem/gate_and.sym
** sch_path: /foss/designs/chipathon_2025/designs/gf180/gate_and/xschem/gate_and.sch
.subckt gate_and B VDD VSS OUT A
*.PININFO OUT:O A:I VDD:B VSS:B B:I
MNB OUTN B NX VSS nfet_03v3 L=0.28u W=1u nf=1 m=4
MPB OUTN B VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
MNA NX A VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=4
MPA OUTN A VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
MIN OUT OUTN VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MIP OUT OUTN VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
.ends


* expanding   symbol:  gf180/gate_inv_L0d5/xschem/gate_inv_L0d5.sym # of pins=4
** sym_path: /foss/designs/chipathon_2025/designs/gf180/gate_inv_L0d5/xschem/gate_inv_L0d5.sym
** sch_path: /foss/designs/chipathon_2025/designs/gf180/gate_inv_L0d5/xschem/gate_inv_L0d5.sch
.subckt gate_inv_L0d5 VDD B A VSS
*.PININFO B:O A:I VDD:B VSS:B
MN B A VSS VSS nfet_03v3 L=0.5u W=1u nf=1 m=2
MP B A VDD VDD pfet_03v3 L=0.5u W=3u nf=1 m=2
.ends

