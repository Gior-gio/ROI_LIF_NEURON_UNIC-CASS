** sch_path: /foss/designs/chipathon_2025/designs/gf180/gate_or/xschem/gate_or.sch
.subckt gate_or B VDD VSS OUT A
*.PININFO OUT:O A:I VDD:B VSS:B B:I
MNB OUTN B VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MPB OUTN B net1 VDD pfet_03v3 L=0.28u W=3u nf=1 m=4
MNA OUTN A VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MPA net1 A VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=4
MIN OUT OUTN VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MIP OUT OUTN VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
MPB1 net1 VDD VDD VDD pfet_03v3 L=0.28u W=3u nf=1 m=2
MNA1 OUTN VSS VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=2
MNA2 VSS VSS VSS VSS nfet_03v3 L=0.28u W=1u nf=1 m=4
.ends
