* Extracted by KLayout with GF180MCU LVS runset on : 19/11/2025 00:59

.SUBCKT spike_generator VSS Ven A Vspk Vrst Vcmp VDD
M$1 \$24 Vcmp VDD VDD pfet_03v3 L=0.28U W=6U AS=3.48P AD=2.505P PS=11.32U
+ PD=7.67U
M$3 \$60 \$24 VDD VDD pfet_03v3 L=0.28U W=12U AS=5.16P AD=5.235P PS=15.44U
+ PD=15.49U
M$7 \$60 VDD VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$8 \$4 Ven \$60 VDD pfet_03v3 L=0.28U W=12U AS=5.16P AD=5.16P PS=15.44U
+ PD=15.44U
M$13 A \$4 VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$15 \$13 \$24 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$17 \$14 \$13 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$19 \$15 \$14 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$21 \$16 \$15 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$23 \$17 \$16 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=3.48P PS=7.72U
+ PD=11.32U
M$25 \$40 \$17 VDD VDD pfet_03v3 L=0.28U W=6U AS=3.48P AD=2.58P PS=11.32U
+ PD=7.72U
M$27 \$40 \$24 VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=3.48P PS=7.72U
+ PD=11.32U
M$29 \$47 \$40 VDD VDD pfet_03v3 L=0.28U W=6U AS=3.48P AD=2.58P PS=11.32U
+ PD=7.72U
M$31 \$31 \$47 VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=2.58P PS=7.72U
+ PD=7.72U
M$33 Vspk \$31 VDD VDD pfet_03v3 L=0.28U W=18U AS=7.74P AD=7.74P PS=23.16U
+ PD=23.16U
M$39 \$32 A VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$41 Vrst \$32 VDD VDD pfet_03v3 L=0.28U W=18U AS=7.74P AD=8.64P PS=23.16U
+ PD=26.76U
M$47 \$24 Vcmp VSS VSS nfet_03v3 L=0.28U W=2U AS=1.16P AD=0.86P PS=5.32U
+ PD=3.72U
M$49 VSS VSS VSS VSS nfet_03v3 L=0.28U W=4U AS=1.72P AD=1.72P PS=7.44U PD=7.44U
M$50 \$4 \$24 VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$54 \$4 VSS VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$55 VSS Ven \$4 VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$59 A \$4 VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$61 \$13 \$24 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$63 \$14 \$13 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$65 \$15 \$14 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$67 \$16 \$15 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$69 \$17 \$16 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$71 \$36 \$17 VSS VSS nfet_03v3 L=0.28U W=4U AS=1.72P AD=1.72P PS=7.44U
+ PD=7.44U
M$72 \$40 \$24 \$36 VSS nfet_03v3 L=0.28U W=4U AS=1.72P AD=1.72P PS=7.44U
+ PD=7.44U
M$79 \$47 \$40 VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U
+ PD=3.72U
M$81 \$31 \$47 VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U
+ PD=3.72U
M$83 Vspk \$31 VSS VSS nfet_03v3 L=0.28U W=6U AS=2.58P AD=2.58P PS=11.16U
+ PD=11.16U
M$89 \$32 A VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$91 Vrst \$32 VSS VSS nfet_03v3 L=0.28U W=6U AS=2.58P AD=2.88P PS=11.16U
+ PD=12.76U
.ENDS spike_generator
