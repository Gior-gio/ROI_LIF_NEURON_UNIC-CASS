* Extracted by KLayout with SG13G2 LVS runset on : 29/01/2026 23:24

.SUBCKT gate_buff_L0d13 VSS VOUT VIN VDD
M$1 VSS VIN \$2 VSS sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$2 VSS \$2 VOUT VSS sg13_lv_nmos L=0.13u W=3u AS=0.72p AD=0.72p PS=5.44u
+ PD=5.44u
M$5 VDD VIN \$2 VDD sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$6 VDD \$2 VOUT VDD sg13_lv_pmos L=0.13u W=6u AS=1.44p AD=1.44p PS=9.44u
+ PD=9.44u
.ENDS gate_buff_L0d13
