* Extracted by KLayout with GF180MCU LVS runset on : 16/11/2025 03:43

.SUBCKT gate_and VSS B A OUT VDD
M$1 \$5 A VDD VDD pfet_03v3 L=0.28U W=6U AS=3.48P AD=2.58P PS=11.32U PD=7.72U
M$3 \$5 B VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=3.48P PS=7.72U PD=11.32U
M$5 OUT \$5 VDD VDD pfet_03v3 L=0.28U W=6U AS=3.48P AD=3.48P PS=11.32U PD=11.32U
M$7 \$4 A VSS VSS nfet_03v3 L=0.28U W=4U AS=2.02P AD=1.72P PS=9.04U PD=7.44U
M$8 \$5 B \$4 VSS nfet_03v3 L=0.28U W=4U AS=1.72P AD=1.72P PS=7.44U PD=7.44U
M$15 OUT \$5 VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=1.16P PS=3.72U PD=5.32U
.ENDS gate_and
