* Extracted by KLayout with GF180MCU LVS runset on : 16/11/2025 06:06

.SUBCKT edge_detector_TOP VSS IN OUT VDD
M$1 OUT \$13 VDD VDD pfet_03v3 L=0.28U W=6U AS=3.48P AD=3.48P PS=11.32U
+ PD=11.32U
M$3 \$13 \$8 VDD VDD pfet_03v3 L=0.28U W=6U AS=3.48P AD=2.58P PS=11.32U PD=7.72U
M$5 \$13 IN VDD VDD pfet_03v3 L=0.28U W=6U AS=2.58P AD=3.48P PS=7.72U PD=11.32U
M$7 \$3 IN VDD VDD pfet_03v3 L=0.5U W=6U AS=3.48P AD=2.58P PS=11.32U PD=7.72U
M$9 \$5 \$3 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$11 \$6 \$5 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$13 \$7 \$6 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=2.58P PS=7.72U PD=7.72U
M$15 \$8 \$7 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.58P AD=3.48P PS=7.72U PD=11.32U
M$17 \$3 IN VSS VSS nfet_03v3 L=0.5U W=2U AS=1.16P AD=0.86P PS=5.32U PD=3.72U
M$19 \$5 \$3 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$21 \$6 \$5 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$23 \$7 \$6 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$25 \$8 \$7 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.86P AD=0.86P PS=3.72U PD=3.72U
M$27 \$14 \$8 VSS VSS nfet_03v3 L=0.28U W=4U AS=1.72P AD=1.72P PS=7.44U PD=7.44U
M$28 \$13 IN \$14 VSS nfet_03v3 L=0.28U W=4U AS=1.72P AD=1.72P PS=7.44U PD=7.44U
M$35 OUT \$13 VSS VSS nfet_03v3 L=0.28U W=2U AS=0.86P AD=1.16P PS=3.72U PD=5.32U
.ENDS edge_detector_TOP
